/*
 Produced by NSL Core(version=20151214), IP ARCH, Inc. Thu Mar 15 10:14:03 2018
 Licensed to :EVALUATION USER
*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module receiver ( m_clock , p_reset );
  input m_clock;
  wire m_clock;
  input p_reset;
  wire p_reset;

endmodule
/*
 Produced by NSL Core(version=20151214), IP ARCH, Inc. Thu Mar 15 10:14:03 2018
 Licensed to :EVALUATION USER
*/
